module game_over_screen (
input px,
input py,

output pixels);



endmodule