module collision_detector(
);

endmodule
