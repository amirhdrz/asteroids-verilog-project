module Rocks(
input [9:0] x,
input [9:0] y,
output [9:0] red, 
output [9:0] green, 
output [9:0] blue,
input clk,
);


endmodule